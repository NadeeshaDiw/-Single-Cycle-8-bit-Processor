//testbench for the ALU module
module testbed;

	//definning signals that are needed to instantiate the ALU module
	reg [7:0] OPERAND1, OPERAND2;
	wire [7:0] ALURESULT;
	reg [2:0] ALUOP;
	
	//set to monitor the values in the signals
	initial begin
		$monitor ($time, " Operand-1 =%d,	Operand-2 =%d,	ALU-OP =%b,	ALU-Result =%d", OPERAND1, OPERAND2, ALUOP, ALURESULT);
	end
	
	//instantiate the ALU module
	alu a1(OPERAND1, OPERAND2, ALURESULT, ALUOP);

	//set values to the signals
	initial
	begin
		$dumpfile("alu.vcd");
		$dumpvars(0, testbed);
	
		OPERAND1 = 8'b0010_0001;
		OPERAND2 = 8'b0100_0011;
		#10 ALUOP = 3'b000;
		#10 ALUOP = 3'b001;
		#10 ALUOP = 3'b010;
		#10 ALUOP = 3'b011;
		#10 ALUOP = 3'b100;
		OPERAND1 = 8'b1010_1111;
		OPERAND2 = 8'b0100_1011;
		#10 ALUOP = 3'b000;
		#10 ALUOP = 3'b001;
		#10 ALUOP = 3'b010;
		#10 ALUOP = 3'b011;
		#10 ALUOP = 3'b100;
	end
	
	//set the simulation life
	initial
	begin
		#100 $finish;	//after 100 units of simulation time, the simulation will end
	end
	
endmodule

//The ALU module implementation
module alu (DATA1, DATA2, RESULT, SELECT);

	//definning input ports
	input [7:0] DATA1, DATA2;
	input [2:0] SELECT;

	//definning output ports
	output reg [7:0] RESULT;
	
	//definning temparary wires to carry the result generated by each functional modules
	wire [7:0] RESULT_FW, RESULT_AD, RESULT_AND, RESULT_OR;
	
	//instantiating the each functional modules
	FORWARD fw (DATA2, RESULT_FW);
	ADD ad (DATA1, DATA2, RESULT_AD);
	AND an (DATA1, DATA2, RESULT_AND);
	OR orr (DATA1, DATA2, RESULT_OR);
	
	//The MUX implementation
	always @(DATA1, DATA2, SELECT)	//sensirive ports for the mux
	begin
		//definning case structure to handle the output of the mux according to the select signal
		case (SELECT)	
			3'b000 :	RESULT = RESULT_FW;		//if SELECT = 0; RESULT will get the output of FORWARD functional unit
			3'b001 :	RESULT = RESULT_AD;		//if SELECT = 1; RESULT will get the output of ADD functional unit
			3'b010 :	RESULT = RESULT_AND;	//if SELECT = 2; RESULT will get the output of AND functional unit
			3'b011 :	RESULT = RESULT_OR;		//if SELECT = 3; RESULT will get the output of OR functional unit
			default :	RESULT = 8'b0000_0000;	//if SELECT > 3; RESULT is set to the zero value
		endcase
	end
	
endmodule

//FORWARD function implementation
module FORWARD (DATA2, RESULT);

	input [7:0] DATA2;		//definning input ports
	output reg [7:0] RESULT;	//definning output ports
	
	//Forward operation happens and result is stored in RESULT net
	always @(DATA2)
	begin
		RESULT = #1 DATA2;		//unit delay assign to 1 time unit
	end

endmodule

//ADD function implementation
module ADD (DATA1, DATA2, RESULT);
	
	input [7:0] DATA1, DATA2;	//definning input ports
	output reg [7:0] RESULT;	//definning output ports
	
	//ADD operation happens and result is stored in RESULT net
	always @(DATA1, DATA2)
	begin
		RESULT = #2 (DATA1 + DATA2);		//unit time delay assign to 2 time unit
	end
	
endmodule

//AND function implementation
module AND(DATA1, DATA2, RESULT);
	
	input [7:0] DATA1, DATA2;	//definning input ports
	output reg [7:0] RESULT;	//definning output ports
	
	//AND operation happens and result is stored in RESULT net
	always @(DATA1, DATA2)
	begin
		RESULT = #1 (DATA1 & DATA2);		//unit time delay assign to 1 time unit
	end
	
endmodule

//OR function implementation
module OR (DATA1, DATA2, RESULT);

	input [7:0] DATA1, DATA2;	//definning input ports
	output reg [7:0] RESULT;	//definning output ports
	
	//OR operation happen result is stored in RESULT net
	always @(DATA1, DATA2)
	begin
		RESULT = #1 (DATA1 | DATA2);		//unit time delay assign to 1 time unit
	end

endmodule
